module branch_comp(
    input[31:0] data_in_A,
    input[31:0] data_in_B,
    input brun_sel,
    output reg br_eq,
    output reg br_lt
);
always @( * ) begin
    case(brun_sel)
    1'b0:begin
        br_eq = ($signed(data_in_A) == $signed(data_in_B))? 1:0;
        br_lt = ($signed(data_in_A) < $signed(data_in_B))? 1:0;
    end
    1'b1:begin
        br_eq = ($unsigned(data_in_A) == $unsigned(data_in_B))? 1:0;
        br_lt = ($unsigned(data_in_A) < $unsigned(data_in_B))? 1:0;
    end
    endcase
end
endmodule